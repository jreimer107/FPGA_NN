module Decoder_11_2048(in, out);
	input [11:0] in;
	output [2048:0] out;

	wire A, B, C, D, E, F, G, H, I, J, K;

	assign out[000] = ~A & ~B & ~C & ~D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[001] = ~A & ~B & ~C & ~D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[002] = ~A & ~B & ~C & ~D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[003] = ~A & ~B & ~C & ~D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[004] = ~A & ~B & ~C & ~D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[005] = ~A & ~B & ~C & ~D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[006] = ~A & ~B & ~C & ~D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[007] = ~A & ~B & ~C & ~D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[008] = ~A & ~B & ~C & ~D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[009] = ~A & ~B & ~C & ~D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[010] = ~A & ~B & ~C & ~D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[011] = ~A & ~B & ~C & ~D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[012] = ~A & ~B & ~C & ~D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[013] = ~A & ~B & ~C & ~D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[014] = ~A & ~B & ~C & ~D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[015] = ~A & ~B & ~C & ~D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[016] = ~A & ~B & ~C & ~D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[017] = ~A & ~B & ~C & ~D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[018] = ~A & ~B & ~C & ~D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[019] = ~A & ~B & ~C & ~D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[020] = ~A & ~B & ~C & ~D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[021] = ~A & ~B & ~C & ~D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[022] = ~A & ~B & ~C & ~D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[023] = ~A & ~B & ~C & ~D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[024] = ~A & ~B & ~C & ~D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[025] = ~A & ~B & ~C & ~D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[026] = ~A & ~B & ~C & ~D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[027] = ~A & ~B & ~C & ~D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[028] = ~A & ~B & ~C & ~D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[029] = ~A & ~B & ~C & ~D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[030] = ~A & ~B & ~C & ~D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[031] = ~A & ~B & ~C & ~D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[032] = ~A & ~B & ~C & ~D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[033] = ~A & ~B & ~C & ~D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[034] = ~A & ~B & ~C & ~D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[035] = ~A & ~B & ~C & ~D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[036] = ~A & ~B & ~C & ~D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[037] = ~A & ~B & ~C & ~D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[038] = ~A & ~B & ~C & ~D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[039] = ~A & ~B & ~C & ~D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[040] = ~A & ~B & ~C & ~D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[041] = ~A & ~B & ~C & ~D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[042] = ~A & ~B & ~C & ~D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[043] = ~A & ~B & ~C & ~D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[044] = ~A & ~B & ~C & ~D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[045] = ~A & ~B & ~C & ~D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[046] = ~A & ~B & ~C & ~D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[047] = ~A & ~B & ~C & ~D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[048] = ~A & ~B & ~C & ~D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[049] = ~A & ~B & ~C & ~D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[050] = ~A & ~B & ~C & ~D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[051] = ~A & ~B & ~C & ~D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[052] = ~A & ~B & ~C & ~D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[053] = ~A & ~B & ~C & ~D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[054] = ~A & ~B & ~C & ~D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[055] = ~A & ~B & ~C & ~D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[056] = ~A & ~B & ~C & ~D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[057] = ~A & ~B & ~C & ~D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[058] = ~A & ~B & ~C & ~D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[059] = ~A & ~B & ~C & ~D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[060] = ~A & ~B & ~C & ~D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[061] = ~A & ~B & ~C & ~D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[062] = ~A & ~B & ~C & ~D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[063] = ~A & ~B & ~C & ~D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[064] = ~A & ~B & ~C & ~D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[065] = ~A & ~B & ~C & ~D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[066] = ~A & ~B & ~C & ~D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[067] = ~A & ~B & ~C & ~D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[068] = ~A & ~B & ~C & ~D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[069] = ~A & ~B & ~C & ~D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[070] = ~A & ~B & ~C & ~D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[071] = ~A & ~B & ~C & ~D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[072] = ~A & ~B & ~C & ~D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[073] = ~A & ~B & ~C & ~D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[074] = ~A & ~B & ~C & ~D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[075] = ~A & ~B & ~C & ~D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[076] = ~A & ~B & ~C & ~D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[077] = ~A & ~B & ~C & ~D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[078] = ~A & ~B & ~C & ~D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[079] = ~A & ~B & ~C & ~D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[080] = ~A & ~B & ~C & ~D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[081] = ~A & ~B & ~C & ~D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[082] = ~A & ~B & ~C & ~D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[083] = ~A & ~B & ~C & ~D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[084] = ~A & ~B & ~C & ~D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[085] = ~A & ~B & ~C & ~D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[086] = ~A & ~B & ~C & ~D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[087] = ~A & ~B & ~C & ~D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[088] = ~A & ~B & ~C & ~D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[089] = ~A & ~B & ~C & ~D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[090] = ~A & ~B & ~C & ~D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[091] = ~A & ~B & ~C & ~D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[092] = ~A & ~B & ~C & ~D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[093] = ~A & ~B & ~C & ~D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[094] = ~A & ~B & ~C & ~D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[095] = ~A & ~B & ~C & ~D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[096] = ~A & ~B & ~C & ~D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[097] = ~A & ~B & ~C & ~D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[098] = ~A & ~B & ~C & ~D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[099] = ~A & ~B & ~C & ~D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[100] = ~A & ~B & ~C & ~D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[101] = ~A & ~B & ~C & ~D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[102] = ~A & ~B & ~C & ~D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[103] = ~A & ~B & ~C & ~D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[104] = ~A & ~B & ~C & ~D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[105] = ~A & ~B & ~C & ~D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[106] = ~A & ~B & ~C & ~D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[107] = ~A & ~B & ~C & ~D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[108] = ~A & ~B & ~C & ~D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[109] = ~A & ~B & ~C & ~D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[110] = ~A & ~B & ~C & ~D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[111] = ~A & ~B & ~C & ~D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[112] = ~A & ~B & ~C & ~D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[113] = ~A & ~B & ~C & ~D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[114] = ~A & ~B & ~C & ~D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[115] = ~A & ~B & ~C & ~D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[116] = ~A & ~B & ~C & ~D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[117] = ~A & ~B & ~C & ~D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[118] = ~A & ~B & ~C & ~D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[119] = ~A & ~B & ~C & ~D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[120] = ~A & ~B & ~C & ~D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[121] = ~A & ~B & ~C & ~D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[122] = ~A & ~B & ~C & ~D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[123] = ~A & ~B & ~C & ~D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[124] = ~A & ~B & ~C & ~D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[125] = ~A & ~B & ~C & ~D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[126] = ~A & ~B & ~C & ~D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[127] = ~A & ~B & ~C & ~D &  E &  F &  G &  H &  I &  J &  K;
	assign out[128] = ~A & ~B & ~C &  D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[129] = ~A & ~B & ~C &  D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[130] = ~A & ~B & ~C &  D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[131] = ~A & ~B & ~C &  D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[132] = ~A & ~B & ~C &  D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[133] = ~A & ~B & ~C &  D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[134] = ~A & ~B & ~C &  D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[135] = ~A & ~B & ~C &  D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[136] = ~A & ~B & ~C &  D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[137] = ~A & ~B & ~C &  D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[138] = ~A & ~B & ~C &  D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[139] = ~A & ~B & ~C &  D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[140] = ~A & ~B & ~C &  D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[141] = ~A & ~B & ~C &  D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[142] = ~A & ~B & ~C &  D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[143] = ~A & ~B & ~C &  D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[144] = ~A & ~B & ~C &  D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[145] = ~A & ~B & ~C &  D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[146] = ~A & ~B & ~C &  D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[147] = ~A & ~B & ~C &  D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[148] = ~A & ~B & ~C &  D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[149] = ~A & ~B & ~C &  D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[150] = ~A & ~B & ~C &  D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[151] = ~A & ~B & ~C &  D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[152] = ~A & ~B & ~C &  D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[153] = ~A & ~B & ~C &  D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[154] = ~A & ~B & ~C &  D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[155] = ~A & ~B & ~C &  D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[156] = ~A & ~B & ~C &  D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[157] = ~A & ~B & ~C &  D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[158] = ~A & ~B & ~C &  D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[159] = ~A & ~B & ~C &  D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[160] = ~A & ~B & ~C &  D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[161] = ~A & ~B & ~C &  D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[162] = ~A & ~B & ~C &  D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[163] = ~A & ~B & ~C &  D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[164] = ~A & ~B & ~C &  D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[165] = ~A & ~B & ~C &  D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[166] = ~A & ~B & ~C &  D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[167] = ~A & ~B & ~C &  D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[168] = ~A & ~B & ~C &  D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[169] = ~A & ~B & ~C &  D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[170] = ~A & ~B & ~C &  D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[171] = ~A & ~B & ~C &  D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[172] = ~A & ~B & ~C &  D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[173] = ~A & ~B & ~C &  D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[174] = ~A & ~B & ~C &  D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[175] = ~A & ~B & ~C &  D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[176] = ~A & ~B & ~C &  D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[177] = ~A & ~B & ~C &  D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[178] = ~A & ~B & ~C &  D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[179] = ~A & ~B & ~C &  D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[180] = ~A & ~B & ~C &  D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[181] = ~A & ~B & ~C &  D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[182] = ~A & ~B & ~C &  D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[183] = ~A & ~B & ~C &  D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[184] = ~A & ~B & ~C &  D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[185] = ~A & ~B & ~C &  D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[186] = ~A & ~B & ~C &  D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[187] = ~A & ~B & ~C &  D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[188] = ~A & ~B & ~C &  D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[189] = ~A & ~B & ~C &  D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[190] = ~A & ~B & ~C &  D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[191] = ~A & ~B & ~C &  D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[192] = ~A & ~B & ~C &  D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[193] = ~A & ~B & ~C &  D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[194] = ~A & ~B & ~C &  D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[195] = ~A & ~B & ~C &  D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[196] = ~A & ~B & ~C &  D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[197] = ~A & ~B & ~C &  D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[198] = ~A & ~B & ~C &  D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[199] = ~A & ~B & ~C &  D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[200] = ~A & ~B & ~C &  D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[201] = ~A & ~B & ~C &  D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[202] = ~A & ~B & ~C &  D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[203] = ~A & ~B & ~C &  D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[204] = ~A & ~B & ~C &  D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[205] = ~A & ~B & ~C &  D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[206] = ~A & ~B & ~C &  D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[207] = ~A & ~B & ~C &  D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[208] = ~A & ~B & ~C &  D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[209] = ~A & ~B & ~C &  D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[210] = ~A & ~B & ~C &  D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[211] = ~A & ~B & ~C &  D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[212] = ~A & ~B & ~C &  D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[213] = ~A & ~B & ~C &  D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[214] = ~A & ~B & ~C &  D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[215] = ~A & ~B & ~C &  D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[216] = ~A & ~B & ~C &  D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[217] = ~A & ~B & ~C &  D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[218] = ~A & ~B & ~C &  D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[219] = ~A & ~B & ~C &  D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[220] = ~A & ~B & ~C &  D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[221] = ~A & ~B & ~C &  D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[222] = ~A & ~B & ~C &  D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[223] = ~A & ~B & ~C &  D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[224] = ~A & ~B & ~C &  D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[225] = ~A & ~B & ~C &  D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[226] = ~A & ~B & ~C &  D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[227] = ~A & ~B & ~C &  D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[228] = ~A & ~B & ~C &  D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[229] = ~A & ~B & ~C &  D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[230] = ~A & ~B & ~C &  D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[231] = ~A & ~B & ~C &  D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[232] = ~A & ~B & ~C &  D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[233] = ~A & ~B & ~C &  D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[234] = ~A & ~B & ~C &  D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[235] = ~A & ~B & ~C &  D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[236] = ~A & ~B & ~C &  D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[237] = ~A & ~B & ~C &  D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[238] = ~A & ~B & ~C &  D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[239] = ~A & ~B & ~C &  D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[240] = ~A & ~B & ~C &  D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[241] = ~A & ~B & ~C &  D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[242] = ~A & ~B & ~C &  D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[243] = ~A & ~B & ~C &  D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[244] = ~A & ~B & ~C &  D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[245] = ~A & ~B & ~C &  D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[246] = ~A & ~B & ~C &  D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[247] = ~A & ~B & ~C &  D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[248] = ~A & ~B & ~C &  D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[249] = ~A & ~B & ~C &  D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[250] = ~A & ~B & ~C &  D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[251] = ~A & ~B & ~C &  D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[252] = ~A & ~B & ~C &  D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[253] = ~A & ~B & ~C &  D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[254] = ~A & ~B & ~C &  D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[255] = ~A & ~B & ~C &  D &  E &  F &  G &  H &  I &  J &  K;
	assign out[256] = ~A & ~B &  C & ~D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[257] = ~A & ~B &  C & ~D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[258] = ~A & ~B &  C & ~D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[259] = ~A & ~B &  C & ~D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[260] = ~A & ~B &  C & ~D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[261] = ~A & ~B &  C & ~D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[262] = ~A & ~B &  C & ~D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[263] = ~A & ~B &  C & ~D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[264] = ~A & ~B &  C & ~D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[265] = ~A & ~B &  C & ~D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[266] = ~A & ~B &  C & ~D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[267] = ~A & ~B &  C & ~D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[268] = ~A & ~B &  C & ~D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[269] = ~A & ~B &  C & ~D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[270] = ~A & ~B &  C & ~D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[271] = ~A & ~B &  C & ~D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[272] = ~A & ~B &  C & ~D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[273] = ~A & ~B &  C & ~D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[274] = ~A & ~B &  C & ~D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[275] = ~A & ~B &  C & ~D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[276] = ~A & ~B &  C & ~D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[277] = ~A & ~B &  C & ~D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[278] = ~A & ~B &  C & ~D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[279] = ~A & ~B &  C & ~D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[280] = ~A & ~B &  C & ~D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[281] = ~A & ~B &  C & ~D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[282] = ~A & ~B &  C & ~D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[283] = ~A & ~B &  C & ~D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[284] = ~A & ~B &  C & ~D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[285] = ~A & ~B &  C & ~D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[286] = ~A & ~B &  C & ~D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[287] = ~A & ~B &  C & ~D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[288] = ~A & ~B &  C & ~D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[289] = ~A & ~B &  C & ~D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[290] = ~A & ~B &  C & ~D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[291] = ~A & ~B &  C & ~D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[292] = ~A & ~B &  C & ~D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[293] = ~A & ~B &  C & ~D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[294] = ~A & ~B &  C & ~D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[295] = ~A & ~B &  C & ~D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[296] = ~A & ~B &  C & ~D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[297] = ~A & ~B &  C & ~D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[298] = ~A & ~B &  C & ~D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[299] = ~A & ~B &  C & ~D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[300] = ~A & ~B &  C & ~D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[301] = ~A & ~B &  C & ~D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[302] = ~A & ~B &  C & ~D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[303] = ~A & ~B &  C & ~D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[304] = ~A & ~B &  C & ~D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[305] = ~A & ~B &  C & ~D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[306] = ~A & ~B &  C & ~D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[307] = ~A & ~B &  C & ~D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[308] = ~A & ~B &  C & ~D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[309] = ~A & ~B &  C & ~D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[310] = ~A & ~B &  C & ~D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[311] = ~A & ~B &  C & ~D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[312] = ~A & ~B &  C & ~D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[313] = ~A & ~B &  C & ~D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[314] = ~A & ~B &  C & ~D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[315] = ~A & ~B &  C & ~D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[316] = ~A & ~B &  C & ~D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[317] = ~A & ~B &  C & ~D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[318] = ~A & ~B &  C & ~D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[319] = ~A & ~B &  C & ~D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[320] = ~A & ~B &  C & ~D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[321] = ~A & ~B &  C & ~D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[322] = ~A & ~B &  C & ~D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[323] = ~A & ~B &  C & ~D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[324] = ~A & ~B &  C & ~D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[325] = ~A & ~B &  C & ~D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[326] = ~A & ~B &  C & ~D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[327] = ~A & ~B &  C & ~D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[328] = ~A & ~B &  C & ~D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[329] = ~A & ~B &  C & ~D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[330] = ~A & ~B &  C & ~D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[331] = ~A & ~B &  C & ~D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[332] = ~A & ~B &  C & ~D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[333] = ~A & ~B &  C & ~D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[334] = ~A & ~B &  C & ~D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[335] = ~A & ~B &  C & ~D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[336] = ~A & ~B &  C & ~D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[337] = ~A & ~B &  C & ~D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[338] = ~A & ~B &  C & ~D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[339] = ~A & ~B &  C & ~D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[340] = ~A & ~B &  C & ~D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[341] = ~A & ~B &  C & ~D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[342] = ~A & ~B &  C & ~D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[343] = ~A & ~B &  C & ~D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[344] = ~A & ~B &  C & ~D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[345] = ~A & ~B &  C & ~D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[346] = ~A & ~B &  C & ~D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[347] = ~A & ~B &  C & ~D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[348] = ~A & ~B &  C & ~D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[349] = ~A & ~B &  C & ~D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[350] = ~A & ~B &  C & ~D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[351] = ~A & ~B &  C & ~D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[352] = ~A & ~B &  C & ~D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[353] = ~A & ~B &  C & ~D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[354] = ~A & ~B &  C & ~D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[355] = ~A & ~B &  C & ~D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[356] = ~A & ~B &  C & ~D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[357] = ~A & ~B &  C & ~D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[358] = ~A & ~B &  C & ~D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[359] = ~A & ~B &  C & ~D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[360] = ~A & ~B &  C & ~D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[361] = ~A & ~B &  C & ~D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[362] = ~A & ~B &  C & ~D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[363] = ~A & ~B &  C & ~D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[364] = ~A & ~B &  C & ~D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[365] = ~A & ~B &  C & ~D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[366] = ~A & ~B &  C & ~D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[367] = ~A & ~B &  C & ~D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[368] = ~A & ~B &  C & ~D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[369] = ~A & ~B &  C & ~D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[370] = ~A & ~B &  C & ~D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[371] = ~A & ~B &  C & ~D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[372] = ~A & ~B &  C & ~D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[373] = ~A & ~B &  C & ~D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[374] = ~A & ~B &  C & ~D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[375] = ~A & ~B &  C & ~D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[376] = ~A & ~B &  C & ~D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[377] = ~A & ~B &  C & ~D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[378] = ~A & ~B &  C & ~D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[379] = ~A & ~B &  C & ~D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[380] = ~A & ~B &  C & ~D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[381] = ~A & ~B &  C & ~D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[382] = ~A & ~B &  C & ~D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[383] = ~A & ~B &  C & ~D &  E &  F &  G &  H &  I &  J &  K;
	assign out[384] = ~A & ~B &  C &  D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[385] = ~A & ~B &  C &  D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[386] = ~A & ~B &  C &  D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[387] = ~A & ~B &  C &  D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[388] = ~A & ~B &  C &  D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[389] = ~A & ~B &  C &  D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[390] = ~A & ~B &  C &  D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[391] = ~A & ~B &  C &  D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[392] = ~A & ~B &  C &  D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[393] = ~A & ~B &  C &  D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[394] = ~A & ~B &  C &  D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[395] = ~A & ~B &  C &  D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[396] = ~A & ~B &  C &  D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[397] = ~A & ~B &  C &  D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[398] = ~A & ~B &  C &  D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[399] = ~A & ~B &  C &  D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[400] = ~A & ~B &  C &  D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[401] = ~A & ~B &  C &  D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[402] = ~A & ~B &  C &  D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[403] = ~A & ~B &  C &  D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[404] = ~A & ~B &  C &  D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[405] = ~A & ~B &  C &  D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[406] = ~A & ~B &  C &  D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[407] = ~A & ~B &  C &  D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[408] = ~A & ~B &  C &  D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[409] = ~A & ~B &  C &  D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[410] = ~A & ~B &  C &  D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[411] = ~A & ~B &  C &  D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[412] = ~A & ~B &  C &  D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[413] = ~A & ~B &  C &  D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[414] = ~A & ~B &  C &  D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[415] = ~A & ~B &  C &  D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[416] = ~A & ~B &  C &  D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[417] = ~A & ~B &  C &  D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[418] = ~A & ~B &  C &  D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[419] = ~A & ~B &  C &  D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[420] = ~A & ~B &  C &  D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[421] = ~A & ~B &  C &  D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[422] = ~A & ~B &  C &  D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[423] = ~A & ~B &  C &  D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[424] = ~A & ~B &  C &  D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[425] = ~A & ~B &  C &  D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[426] = ~A & ~B &  C &  D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[427] = ~A & ~B &  C &  D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[428] = ~A & ~B &  C &  D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[429] = ~A & ~B &  C &  D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[430] = ~A & ~B &  C &  D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[431] = ~A & ~B &  C &  D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[432] = ~A & ~B &  C &  D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[433] = ~A & ~B &  C &  D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[434] = ~A & ~B &  C &  D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[435] = ~A & ~B &  C &  D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[436] = ~A & ~B &  C &  D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[437] = ~A & ~B &  C &  D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[438] = ~A & ~B &  C &  D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[439] = ~A & ~B &  C &  D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[440] = ~A & ~B &  C &  D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[441] = ~A & ~B &  C &  D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[442] = ~A & ~B &  C &  D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[443] = ~A & ~B &  C &  D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[444] = ~A & ~B &  C &  D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[445] = ~A & ~B &  C &  D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[446] = ~A & ~B &  C &  D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[447] = ~A & ~B &  C &  D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[448] = ~A & ~B &  C &  D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[449] = ~A & ~B &  C &  D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[450] = ~A & ~B &  C &  D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[451] = ~A & ~B &  C &  D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[452] = ~A & ~B &  C &  D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[453] = ~A & ~B &  C &  D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[454] = ~A & ~B &  C &  D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[455] = ~A & ~B &  C &  D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[456] = ~A & ~B &  C &  D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[457] = ~A & ~B &  C &  D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[458] = ~A & ~B &  C &  D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[459] = ~A & ~B &  C &  D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[460] = ~A & ~B &  C &  D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[461] = ~A & ~B &  C &  D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[462] = ~A & ~B &  C &  D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[463] = ~A & ~B &  C &  D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[464] = ~A & ~B &  C &  D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[465] = ~A & ~B &  C &  D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[466] = ~A & ~B &  C &  D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[467] = ~A & ~B &  C &  D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[468] = ~A & ~B &  C &  D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[469] = ~A & ~B &  C &  D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[470] = ~A & ~B &  C &  D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[471] = ~A & ~B &  C &  D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[472] = ~A & ~B &  C &  D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[473] = ~A & ~B &  C &  D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[474] = ~A & ~B &  C &  D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[475] = ~A & ~B &  C &  D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[476] = ~A & ~B &  C &  D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[477] = ~A & ~B &  C &  D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[478] = ~A & ~B &  C &  D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[479] = ~A & ~B &  C &  D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[480] = ~A & ~B &  C &  D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[481] = ~A & ~B &  C &  D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[482] = ~A & ~B &  C &  D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[483] = ~A & ~B &  C &  D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[484] = ~A & ~B &  C &  D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[485] = ~A & ~B &  C &  D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[486] = ~A & ~B &  C &  D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[487] = ~A & ~B &  C &  D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[488] = ~A & ~B &  C &  D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[489] = ~A & ~B &  C &  D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[490] = ~A & ~B &  C &  D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[491] = ~A & ~B &  C &  D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[492] = ~A & ~B &  C &  D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[493] = ~A & ~B &  C &  D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[494] = ~A & ~B &  C &  D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[495] = ~A & ~B &  C &  D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[496] = ~A & ~B &  C &  D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[497] = ~A & ~B &  C &  D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[498] = ~A & ~B &  C &  D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[499] = ~A & ~B &  C &  D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[500] = ~A & ~B &  C &  D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[501] = ~A & ~B &  C &  D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[502] = ~A & ~B &  C &  D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[503] = ~A & ~B &  C &  D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[504] = ~A & ~B &  C &  D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[505] = ~A & ~B &  C &  D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[506] = ~A & ~B &  C &  D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[507] = ~A & ~B &  C &  D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[508] = ~A & ~B &  C &  D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[509] = ~A & ~B &  C &  D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[510] = ~A & ~B &  C &  D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[511] = ~A & ~B &  C &  D &  E &  F &  G &  H &  I &  J &  K;
	assign out[512] = ~A &  B & ~C & ~D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[513] = ~A &  B & ~C & ~D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[514] = ~A &  B & ~C & ~D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[515] = ~A &  B & ~C & ~D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[516] = ~A &  B & ~C & ~D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[517] = ~A &  B & ~C & ~D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[518] = ~A &  B & ~C & ~D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[519] = ~A &  B & ~C & ~D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[520] = ~A &  B & ~C & ~D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[521] = ~A &  B & ~C & ~D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[522] = ~A &  B & ~C & ~D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[523] = ~A &  B & ~C & ~D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[524] = ~A &  B & ~C & ~D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[525] = ~A &  B & ~C & ~D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[526] = ~A &  B & ~C & ~D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[527] = ~A &  B & ~C & ~D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[528] = ~A &  B & ~C & ~D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[529] = ~A &  B & ~C & ~D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[530] = ~A &  B & ~C & ~D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[531] = ~A &  B & ~C & ~D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[532] = ~A &  B & ~C & ~D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[533] = ~A &  B & ~C & ~D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[534] = ~A &  B & ~C & ~D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[535] = ~A &  B & ~C & ~D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[536] = ~A &  B & ~C & ~D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[537] = ~A &  B & ~C & ~D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[538] = ~A &  B & ~C & ~D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[539] = ~A &  B & ~C & ~D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[540] = ~A &  B & ~C & ~D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[541] = ~A &  B & ~C & ~D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[542] = ~A &  B & ~C & ~D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[543] = ~A &  B & ~C & ~D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[544] = ~A &  B & ~C & ~D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[545] = ~A &  B & ~C & ~D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[546] = ~A &  B & ~C & ~D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[547] = ~A &  B & ~C & ~D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[548] = ~A &  B & ~C & ~D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[549] = ~A &  B & ~C & ~D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[550] = ~A &  B & ~C & ~D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[551] = ~A &  B & ~C & ~D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[552] = ~A &  B & ~C & ~D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[553] = ~A &  B & ~C & ~D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[554] = ~A &  B & ~C & ~D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[555] = ~A &  B & ~C & ~D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[556] = ~A &  B & ~C & ~D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[557] = ~A &  B & ~C & ~D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[558] = ~A &  B & ~C & ~D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[559] = ~A &  B & ~C & ~D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[560] = ~A &  B & ~C & ~D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[561] = ~A &  B & ~C & ~D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[562] = ~A &  B & ~C & ~D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[563] = ~A &  B & ~C & ~D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[564] = ~A &  B & ~C & ~D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[565] = ~A &  B & ~C & ~D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[566] = ~A &  B & ~C & ~D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[567] = ~A &  B & ~C & ~D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[568] = ~A &  B & ~C & ~D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[569] = ~A &  B & ~C & ~D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[570] = ~A &  B & ~C & ~D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[571] = ~A &  B & ~C & ~D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[572] = ~A &  B & ~C & ~D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[573] = ~A &  B & ~C & ~D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[574] = ~A &  B & ~C & ~D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[575] = ~A &  B & ~C & ~D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[576] = ~A &  B & ~C & ~D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[577] = ~A &  B & ~C & ~D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[578] = ~A &  B & ~C & ~D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[579] = ~A &  B & ~C & ~D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[580] = ~A &  B & ~C & ~D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[581] = ~A &  B & ~C & ~D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[582] = ~A &  B & ~C & ~D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[583] = ~A &  B & ~C & ~D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[584] = ~A &  B & ~C & ~D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[585] = ~A &  B & ~C & ~D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[586] = ~A &  B & ~C & ~D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[587] = ~A &  B & ~C & ~D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[588] = ~A &  B & ~C & ~D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[589] = ~A &  B & ~C & ~D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[590] = ~A &  B & ~C & ~D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[591] = ~A &  B & ~C & ~D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[592] = ~A &  B & ~C & ~D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[593] = ~A &  B & ~C & ~D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[594] = ~A &  B & ~C & ~D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[595] = ~A &  B & ~C & ~D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[596] = ~A &  B & ~C & ~D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[597] = ~A &  B & ~C & ~D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[598] = ~A &  B & ~C & ~D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[599] = ~A &  B & ~C & ~D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[600] = ~A &  B & ~C & ~D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[601] = ~A &  B & ~C & ~D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[602] = ~A &  B & ~C & ~D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[603] = ~A &  B & ~C & ~D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[604] = ~A &  B & ~C & ~D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[605] = ~A &  B & ~C & ~D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[606] = ~A &  B & ~C & ~D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[607] = ~A &  B & ~C & ~D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[608] = ~A &  B & ~C & ~D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[609] = ~A &  B & ~C & ~D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[610] = ~A &  B & ~C & ~D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[611] = ~A &  B & ~C & ~D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[612] = ~A &  B & ~C & ~D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[613] = ~A &  B & ~C & ~D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[614] = ~A &  B & ~C & ~D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[615] = ~A &  B & ~C & ~D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[616] = ~A &  B & ~C & ~D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[617] = ~A &  B & ~C & ~D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[618] = ~A &  B & ~C & ~D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[619] = ~A &  B & ~C & ~D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[620] = ~A &  B & ~C & ~D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[621] = ~A &  B & ~C & ~D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[622] = ~A &  B & ~C & ~D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[623] = ~A &  B & ~C & ~D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[624] = ~A &  B & ~C & ~D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[625] = ~A &  B & ~C & ~D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[626] = ~A &  B & ~C & ~D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[627] = ~A &  B & ~C & ~D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[628] = ~A &  B & ~C & ~D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[629] = ~A &  B & ~C & ~D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[630] = ~A &  B & ~C & ~D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[631] = ~A &  B & ~C & ~D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[632] = ~A &  B & ~C & ~D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[633] = ~A &  B & ~C & ~D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[634] = ~A &  B & ~C & ~D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[635] = ~A &  B & ~C & ~D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[636] = ~A &  B & ~C & ~D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[637] = ~A &  B & ~C & ~D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[638] = ~A &  B & ~C & ~D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[639] = ~A &  B & ~C & ~D &  E &  F &  G &  H &  I &  J &  K;
	assign out[640] = ~A &  B & ~C &  D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[641] = ~A &  B & ~C &  D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[642] = ~A &  B & ~C &  D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[643] = ~A &  B & ~C &  D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[644] = ~A &  B & ~C &  D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[645] = ~A &  B & ~C &  D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[646] = ~A &  B & ~C &  D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[647] = ~A &  B & ~C &  D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[648] = ~A &  B & ~C &  D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[649] = ~A &  B & ~C &  D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[650] = ~A &  B & ~C &  D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[651] = ~A &  B & ~C &  D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[652] = ~A &  B & ~C &  D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[653] = ~A &  B & ~C &  D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[654] = ~A &  B & ~C &  D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[655] = ~A &  B & ~C &  D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[656] = ~A &  B & ~C &  D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[657] = ~A &  B & ~C &  D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[658] = ~A &  B & ~C &  D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[659] = ~A &  B & ~C &  D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[660] = ~A &  B & ~C &  D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[661] = ~A &  B & ~C &  D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[662] = ~A &  B & ~C &  D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[663] = ~A &  B & ~C &  D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[664] = ~A &  B & ~C &  D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[665] = ~A &  B & ~C &  D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[666] = ~A &  B & ~C &  D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[667] = ~A &  B & ~C &  D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[668] = ~A &  B & ~C &  D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[669] = ~A &  B & ~C &  D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[670] = ~A &  B & ~C &  D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[671] = ~A &  B & ~C &  D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[672] = ~A &  B & ~C &  D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[673] = ~A &  B & ~C &  D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[674] = ~A &  B & ~C &  D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[675] = ~A &  B & ~C &  D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[676] = ~A &  B & ~C &  D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[677] = ~A &  B & ~C &  D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[678] = ~A &  B & ~C &  D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[679] = ~A &  B & ~C &  D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[680] = ~A &  B & ~C &  D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[681] = ~A &  B & ~C &  D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[682] = ~A &  B & ~C &  D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[683] = ~A &  B & ~C &  D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[684] = ~A &  B & ~C &  D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[685] = ~A &  B & ~C &  D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[686] = ~A &  B & ~C &  D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[687] = ~A &  B & ~C &  D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[688] = ~A &  B & ~C &  D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[689] = ~A &  B & ~C &  D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[690] = ~A &  B & ~C &  D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[691] = ~A &  B & ~C &  D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[692] = ~A &  B & ~C &  D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[693] = ~A &  B & ~C &  D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[694] = ~A &  B & ~C &  D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[695] = ~A &  B & ~C &  D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[696] = ~A &  B & ~C &  D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[697] = ~A &  B & ~C &  D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[698] = ~A &  B & ~C &  D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[699] = ~A &  B & ~C &  D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[700] = ~A &  B & ~C &  D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[701] = ~A &  B & ~C &  D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[702] = ~A &  B & ~C &  D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[703] = ~A &  B & ~C &  D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[704] = ~A &  B & ~C &  D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[705] = ~A &  B & ~C &  D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[706] = ~A &  B & ~C &  D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[707] = ~A &  B & ~C &  D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[708] = ~A &  B & ~C &  D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[709] = ~A &  B & ~C &  D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[710] = ~A &  B & ~C &  D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[711] = ~A &  B & ~C &  D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[712] = ~A &  B & ~C &  D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[713] = ~A &  B & ~C &  D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[714] = ~A &  B & ~C &  D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[715] = ~A &  B & ~C &  D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[716] = ~A &  B & ~C &  D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[717] = ~A &  B & ~C &  D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[718] = ~A &  B & ~C &  D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[719] = ~A &  B & ~C &  D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[720] = ~A &  B & ~C &  D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[721] = ~A &  B & ~C &  D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[722] = ~A &  B & ~C &  D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[723] = ~A &  B & ~C &  D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[724] = ~A &  B & ~C &  D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[725] = ~A &  B & ~C &  D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[726] = ~A &  B & ~C &  D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[727] = ~A &  B & ~C &  D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[728] = ~A &  B & ~C &  D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[729] = ~A &  B & ~C &  D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[730] = ~A &  B & ~C &  D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[731] = ~A &  B & ~C &  D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[732] = ~A &  B & ~C &  D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[733] = ~A &  B & ~C &  D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[734] = ~A &  B & ~C &  D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[735] = ~A &  B & ~C &  D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[736] = ~A &  B & ~C &  D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[737] = ~A &  B & ~C &  D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[738] = ~A &  B & ~C &  D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[739] = ~A &  B & ~C &  D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[740] = ~A &  B & ~C &  D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[741] = ~A &  B & ~C &  D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[742] = ~A &  B & ~C &  D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[743] = ~A &  B & ~C &  D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[744] = ~A &  B & ~C &  D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[745] = ~A &  B & ~C &  D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[746] = ~A &  B & ~C &  D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[747] = ~A &  B & ~C &  D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[748] = ~A &  B & ~C &  D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[749] = ~A &  B & ~C &  D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[750] = ~A &  B & ~C &  D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[751] = ~A &  B & ~C &  D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[752] = ~A &  B & ~C &  D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[753] = ~A &  B & ~C &  D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[754] = ~A &  B & ~C &  D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[755] = ~A &  B & ~C &  D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[756] = ~A &  B & ~C &  D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[757] = ~A &  B & ~C &  D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[758] = ~A &  B & ~C &  D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[759] = ~A &  B & ~C &  D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[760] = ~A &  B & ~C &  D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[761] = ~A &  B & ~C &  D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[762] = ~A &  B & ~C &  D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[763] = ~A &  B & ~C &  D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[764] = ~A &  B & ~C &  D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[765] = ~A &  B & ~C &  D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[766] = ~A &  B & ~C &  D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[767] = ~A &  B & ~C &  D &  E &  F &  G &  H &  I &  J &  K;
	assign out[768] = ~A &  B &  C & ~D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[769] = ~A &  B &  C & ~D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[770] = ~A &  B &  C & ~D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[771] = ~A &  B &  C & ~D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[772] = ~A &  B &  C & ~D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[773] = ~A &  B &  C & ~D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[774] = ~A &  B &  C & ~D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[775] = ~A &  B &  C & ~D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[776] = ~A &  B &  C & ~D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[777] = ~A &  B &  C & ~D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[778] = ~A &  B &  C & ~D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[779] = ~A &  B &  C & ~D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[780] = ~A &  B &  C & ~D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[781] = ~A &  B &  C & ~D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[782] = ~A &  B &  C & ~D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[783] = ~A &  B &  C & ~D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[784] = ~A &  B &  C & ~D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[785] = ~A &  B &  C & ~D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[786] = ~A &  B &  C & ~D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[787] = ~A &  B &  C & ~D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[788] = ~A &  B &  C & ~D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[789] = ~A &  B &  C & ~D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[790] = ~A &  B &  C & ~D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[791] = ~A &  B &  C & ~D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[792] = ~A &  B &  C & ~D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[793] = ~A &  B &  C & ~D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[794] = ~A &  B &  C & ~D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[795] = ~A &  B &  C & ~D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[796] = ~A &  B &  C & ~D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[797] = ~A &  B &  C & ~D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[798] = ~A &  B &  C & ~D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[799] = ~A &  B &  C & ~D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[800] = ~A &  B &  C & ~D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[801] = ~A &  B &  C & ~D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[802] = ~A &  B &  C & ~D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[803] = ~A &  B &  C & ~D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[804] = ~A &  B &  C & ~D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[805] = ~A &  B &  C & ~D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[806] = ~A &  B &  C & ~D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[807] = ~A &  B &  C & ~D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[808] = ~A &  B &  C & ~D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[809] = ~A &  B &  C & ~D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[810] = ~A &  B &  C & ~D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[811] = ~A &  B &  C & ~D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[812] = ~A &  B &  C & ~D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[813] = ~A &  B &  C & ~D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[814] = ~A &  B &  C & ~D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[815] = ~A &  B &  C & ~D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[816] = ~A &  B &  C & ~D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[817] = ~A &  B &  C & ~D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[818] = ~A &  B &  C & ~D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[819] = ~A &  B &  C & ~D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[820] = ~A &  B &  C & ~D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[821] = ~A &  B &  C & ~D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[822] = ~A &  B &  C & ~D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[823] = ~A &  B &  C & ~D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[824] = ~A &  B &  C & ~D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[825] = ~A &  B &  C & ~D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[826] = ~A &  B &  C & ~D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[827] = ~A &  B &  C & ~D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[828] = ~A &  B &  C & ~D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[829] = ~A &  B &  C & ~D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[830] = ~A &  B &  C & ~D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[831] = ~A &  B &  C & ~D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[832] = ~A &  B &  C & ~D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[833] = ~A &  B &  C & ~D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[834] = ~A &  B &  C & ~D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[835] = ~A &  B &  C & ~D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[836] = ~A &  B &  C & ~D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[837] = ~A &  B &  C & ~D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[838] = ~A &  B &  C & ~D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[839] = ~A &  B &  C & ~D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[840] = ~A &  B &  C & ~D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[841] = ~A &  B &  C & ~D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[842] = ~A &  B &  C & ~D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[843] = ~A &  B &  C & ~D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[844] = ~A &  B &  C & ~D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[845] = ~A &  B &  C & ~D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[846] = ~A &  B &  C & ~D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[847] = ~A &  B &  C & ~D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[848] = ~A &  B &  C & ~D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[849] = ~A &  B &  C & ~D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[850] = ~A &  B &  C & ~D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[851] = ~A &  B &  C & ~D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[852] = ~A &  B &  C & ~D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[853] = ~A &  B &  C & ~D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[854] = ~A &  B &  C & ~D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[855] = ~A &  B &  C & ~D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[856] = ~A &  B &  C & ~D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[857] = ~A &  B &  C & ~D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[858] = ~A &  B &  C & ~D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[859] = ~A &  B &  C & ~D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[860] = ~A &  B &  C & ~D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[861] = ~A &  B &  C & ~D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[862] = ~A &  B &  C & ~D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[863] = ~A &  B &  C & ~D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[864] = ~A &  B &  C & ~D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[865] = ~A &  B &  C & ~D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[866] = ~A &  B &  C & ~D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[867] = ~A &  B &  C & ~D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[868] = ~A &  B &  C & ~D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[869] = ~A &  B &  C & ~D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[870] = ~A &  B &  C & ~D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[871] = ~A &  B &  C & ~D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[872] = ~A &  B &  C & ~D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[873] = ~A &  B &  C & ~D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[874] = ~A &  B &  C & ~D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[875] = ~A &  B &  C & ~D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[876] = ~A &  B &  C & ~D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[877] = ~A &  B &  C & ~D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[878] = ~A &  B &  C & ~D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[879] = ~A &  B &  C & ~D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[880] = ~A &  B &  C & ~D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[881] = ~A &  B &  C & ~D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[882] = ~A &  B &  C & ~D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[883] = ~A &  B &  C & ~D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[884] = ~A &  B &  C & ~D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[885] = ~A &  B &  C & ~D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[886] = ~A &  B &  C & ~D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[887] = ~A &  B &  C & ~D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[888] = ~A &  B &  C & ~D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[889] = ~A &  B &  C & ~D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[890] = ~A &  B &  C & ~D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[891] = ~A &  B &  C & ~D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[892] = ~A &  B &  C & ~D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[893] = ~A &  B &  C & ~D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[894] = ~A &  B &  C & ~D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[895] = ~A &  B &  C & ~D &  E &  F &  G &  H &  I &  J &  K;
	assign out[896] = ~A &  B &  C &  D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[897] = ~A &  B &  C &  D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[898] = ~A &  B &  C &  D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[899] = ~A &  B &  C &  D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[900] = ~A &  B &  C &  D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[901] = ~A &  B &  C &  D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[902] = ~A &  B &  C &  D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[903] = ~A &  B &  C &  D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[904] = ~A &  B &  C &  D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[905] = ~A &  B &  C &  D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[906] = ~A &  B &  C &  D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[907] = ~A &  B &  C &  D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[908] = ~A &  B &  C &  D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[909] = ~A &  B &  C &  D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[910] = ~A &  B &  C &  D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[911] = ~A &  B &  C &  D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[912] = ~A &  B &  C &  D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[913] = ~A &  B &  C &  D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[914] = ~A &  B &  C &  D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[915] = ~A &  B &  C &  D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[916] = ~A &  B &  C &  D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[917] = ~A &  B &  C &  D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[918] = ~A &  B &  C &  D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[919] = ~A &  B &  C &  D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[920] = ~A &  B &  C &  D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[921] = ~A &  B &  C &  D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[922] = ~A &  B &  C &  D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[923] = ~A &  B &  C &  D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[924] = ~A &  B &  C &  D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[925] = ~A &  B &  C &  D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[926] = ~A &  B &  C &  D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[927] = ~A &  B &  C &  D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[928] = ~A &  B &  C &  D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[929] = ~A &  B &  C &  D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[930] = ~A &  B &  C &  D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[931] = ~A &  B &  C &  D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[932] = ~A &  B &  C &  D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[933] = ~A &  B &  C &  D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[934] = ~A &  B &  C &  D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[935] = ~A &  B &  C &  D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[936] = ~A &  B &  C &  D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[937] = ~A &  B &  C &  D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[938] = ~A &  B &  C &  D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[939] = ~A &  B &  C &  D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[940] = ~A &  B &  C &  D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[941] = ~A &  B &  C &  D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[942] = ~A &  B &  C &  D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[943] = ~A &  B &  C &  D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[944] = ~A &  B &  C &  D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[945] = ~A &  B &  C &  D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[946] = ~A &  B &  C &  D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[947] = ~A &  B &  C &  D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[948] = ~A &  B &  C &  D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[949] = ~A &  B &  C &  D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[950] = ~A &  B &  C &  D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[951] = ~A &  B &  C &  D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[952] = ~A &  B &  C &  D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[953] = ~A &  B &  C &  D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[954] = ~A &  B &  C &  D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[955] = ~A &  B &  C &  D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[956] = ~A &  B &  C &  D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[957] = ~A &  B &  C &  D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[958] = ~A &  B &  C &  D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[959] = ~A &  B &  C &  D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[960] = ~A &  B &  C &  D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[961] = ~A &  B &  C &  D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[962] = ~A &  B &  C &  D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[963] = ~A &  B &  C &  D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[964] = ~A &  B &  C &  D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[965] = ~A &  B &  C &  D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[966] = ~A &  B &  C &  D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[967] = ~A &  B &  C &  D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[968] = ~A &  B &  C &  D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[969] = ~A &  B &  C &  D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[970] = ~A &  B &  C &  D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[971] = ~A &  B &  C &  D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[972] = ~A &  B &  C &  D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[973] = ~A &  B &  C &  D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[974] = ~A &  B &  C &  D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[975] = ~A &  B &  C &  D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[976] = ~A &  B &  C &  D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[977] = ~A &  B &  C &  D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[978] = ~A &  B &  C &  D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[979] = ~A &  B &  C &  D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[980] = ~A &  B &  C &  D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[981] = ~A &  B &  C &  D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[982] = ~A &  B &  C &  D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[983] = ~A &  B &  C &  D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[984] = ~A &  B &  C &  D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[985] = ~A &  B &  C &  D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[986] = ~A &  B &  C &  D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[987] = ~A &  B &  C &  D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[988] = ~A &  B &  C &  D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[989] = ~A &  B &  C &  D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[990] = ~A &  B &  C &  D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[991] = ~A &  B &  C &  D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[992] = ~A &  B &  C &  D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[993] = ~A &  B &  C &  D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[994] = ~A &  B &  C &  D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[995] = ~A &  B &  C &  D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[996] = ~A &  B &  C &  D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[997] = ~A &  B &  C &  D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[998] = ~A &  B &  C &  D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[999] = ~A &  B &  C &  D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[1000] = ~A &  B &  C &  D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1001] = ~A &  B &  C &  D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1002] = ~A &  B &  C &  D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1003] = ~A &  B &  C &  D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[1004] = ~A &  B &  C &  D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1005] = ~A &  B &  C &  D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[1006] = ~A &  B &  C &  D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[1007] = ~A &  B &  C &  D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[1008] = ~A &  B &  C &  D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1009] = ~A &  B &  C &  D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1010] = ~A &  B &  C &  D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1011] = ~A &  B &  C &  D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[1012] = ~A &  B &  C &  D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1013] = ~A &  B &  C &  D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[1014] = ~A &  B &  C &  D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[1015] = ~A &  B &  C &  D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[1016] = ~A &  B &  C &  D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1017] = ~A &  B &  C &  D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[1018] = ~A &  B &  C &  D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[1019] = ~A &  B &  C &  D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[1020] = ~A &  B &  C &  D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[1021] = ~A &  B &  C &  D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[1022] = ~A &  B &  C &  D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[1023] = ~A &  B &  C &  D &  E &  F &  G &  H &  I &  J &  K;
	assign out[1024] =  A & ~B & ~C & ~D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1025] =  A & ~B & ~C & ~D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1026] =  A & ~B & ~C & ~D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1027] =  A & ~B & ~C & ~D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1028] =  A & ~B & ~C & ~D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1029] =  A & ~B & ~C & ~D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1030] =  A & ~B & ~C & ~D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1031] =  A & ~B & ~C & ~D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1032] =  A & ~B & ~C & ~D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1033] =  A & ~B & ~C & ~D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1034] =  A & ~B & ~C & ~D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1035] =  A & ~B & ~C & ~D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1036] =  A & ~B & ~C & ~D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1037] =  A & ~B & ~C & ~D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1038] =  A & ~B & ~C & ~D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1039] =  A & ~B & ~C & ~D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[1040] =  A & ~B & ~C & ~D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1041] =  A & ~B & ~C & ~D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1042] =  A & ~B & ~C & ~D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1043] =  A & ~B & ~C & ~D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1044] =  A & ~B & ~C & ~D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1045] =  A & ~B & ~C & ~D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1046] =  A & ~B & ~C & ~D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1047] =  A & ~B & ~C & ~D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[1048] =  A & ~B & ~C & ~D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1049] =  A & ~B & ~C & ~D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1050] =  A & ~B & ~C & ~D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1051] =  A & ~B & ~C & ~D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[1052] =  A & ~B & ~C & ~D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1053] =  A & ~B & ~C & ~D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[1054] =  A & ~B & ~C & ~D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[1055] =  A & ~B & ~C & ~D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[1056] =  A & ~B & ~C & ~D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1057] =  A & ~B & ~C & ~D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1058] =  A & ~B & ~C & ~D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1059] =  A & ~B & ~C & ~D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1060] =  A & ~B & ~C & ~D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1061] =  A & ~B & ~C & ~D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1062] =  A & ~B & ~C & ~D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1063] =  A & ~B & ~C & ~D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[1064] =  A & ~B & ~C & ~D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1065] =  A & ~B & ~C & ~D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1066] =  A & ~B & ~C & ~D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1067] =  A & ~B & ~C & ~D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[1068] =  A & ~B & ~C & ~D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1069] =  A & ~B & ~C & ~D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[1070] =  A & ~B & ~C & ~D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[1071] =  A & ~B & ~C & ~D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[1072] =  A & ~B & ~C & ~D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1073] =  A & ~B & ~C & ~D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1074] =  A & ~B & ~C & ~D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1075] =  A & ~B & ~C & ~D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[1076] =  A & ~B & ~C & ~D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1077] =  A & ~B & ~C & ~D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[1078] =  A & ~B & ~C & ~D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[1079] =  A & ~B & ~C & ~D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[1080] =  A & ~B & ~C & ~D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1081] =  A & ~B & ~C & ~D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[1082] =  A & ~B & ~C & ~D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[1083] =  A & ~B & ~C & ~D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[1084] =  A & ~B & ~C & ~D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[1085] =  A & ~B & ~C & ~D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[1086] =  A & ~B & ~C & ~D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[1087] =  A & ~B & ~C & ~D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[1088] =  A & ~B & ~C & ~D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1089] =  A & ~B & ~C & ~D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1090] =  A & ~B & ~C & ~D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1091] =  A & ~B & ~C & ~D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1092] =  A & ~B & ~C & ~D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1093] =  A & ~B & ~C & ~D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1094] =  A & ~B & ~C & ~D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1095] =  A & ~B & ~C & ~D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1096] =  A & ~B & ~C & ~D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1097] =  A & ~B & ~C & ~D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1098] =  A & ~B & ~C & ~D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1099] =  A & ~B & ~C & ~D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1100] =  A & ~B & ~C & ~D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1101] =  A & ~B & ~C & ~D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1102] =  A & ~B & ~C & ~D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1103] =  A & ~B & ~C & ~D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[1104] =  A & ~B & ~C & ~D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1105] =  A & ~B & ~C & ~D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1106] =  A & ~B & ~C & ~D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1107] =  A & ~B & ~C & ~D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1108] =  A & ~B & ~C & ~D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1109] =  A & ~B & ~C & ~D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1110] =  A & ~B & ~C & ~D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1111] =  A & ~B & ~C & ~D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[1112] =  A & ~B & ~C & ~D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1113] =  A & ~B & ~C & ~D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1114] =  A & ~B & ~C & ~D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1115] =  A & ~B & ~C & ~D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[1116] =  A & ~B & ~C & ~D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1117] =  A & ~B & ~C & ~D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[1118] =  A & ~B & ~C & ~D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[1119] =  A & ~B & ~C & ~D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[1120] =  A & ~B & ~C & ~D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1121] =  A & ~B & ~C & ~D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1122] =  A & ~B & ~C & ~D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1123] =  A & ~B & ~C & ~D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1124] =  A & ~B & ~C & ~D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1125] =  A & ~B & ~C & ~D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1126] =  A & ~B & ~C & ~D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1127] =  A & ~B & ~C & ~D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[1128] =  A & ~B & ~C & ~D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1129] =  A & ~B & ~C & ~D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1130] =  A & ~B & ~C & ~D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1131] =  A & ~B & ~C & ~D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[1132] =  A & ~B & ~C & ~D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1133] =  A & ~B & ~C & ~D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[1134] =  A & ~B & ~C & ~D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[1135] =  A & ~B & ~C & ~D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[1136] =  A & ~B & ~C & ~D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1137] =  A & ~B & ~C & ~D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1138] =  A & ~B & ~C & ~D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1139] =  A & ~B & ~C & ~D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[1140] =  A & ~B & ~C & ~D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1141] =  A & ~B & ~C & ~D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[1142] =  A & ~B & ~C & ~D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[1143] =  A & ~B & ~C & ~D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[1144] =  A & ~B & ~C & ~D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1145] =  A & ~B & ~C & ~D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[1146] =  A & ~B & ~C & ~D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[1147] =  A & ~B & ~C & ~D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[1148] =  A & ~B & ~C & ~D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[1149] =  A & ~B & ~C & ~D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[1150] =  A & ~B & ~C & ~D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[1151] =  A & ~B & ~C & ~D &  E &  F &  G &  H &  I &  J &  K;
	assign out[1152] =  A & ~B & ~C &  D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1153] =  A & ~B & ~C &  D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1154] =  A & ~B & ~C &  D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1155] =  A & ~B & ~C &  D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1156] =  A & ~B & ~C &  D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1157] =  A & ~B & ~C &  D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1158] =  A & ~B & ~C &  D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1159] =  A & ~B & ~C &  D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1160] =  A & ~B & ~C &  D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1161] =  A & ~B & ~C &  D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1162] =  A & ~B & ~C &  D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1163] =  A & ~B & ~C &  D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1164] =  A & ~B & ~C &  D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1165] =  A & ~B & ~C &  D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1166] =  A & ~B & ~C &  D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1167] =  A & ~B & ~C &  D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[1168] =  A & ~B & ~C &  D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1169] =  A & ~B & ~C &  D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1170] =  A & ~B & ~C &  D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1171] =  A & ~B & ~C &  D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1172] =  A & ~B & ~C &  D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1173] =  A & ~B & ~C &  D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1174] =  A & ~B & ~C &  D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1175] =  A & ~B & ~C &  D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[1176] =  A & ~B & ~C &  D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1177] =  A & ~B & ~C &  D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1178] =  A & ~B & ~C &  D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1179] =  A & ~B & ~C &  D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[1180] =  A & ~B & ~C &  D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1181] =  A & ~B & ~C &  D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[1182] =  A & ~B & ~C &  D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[1183] =  A & ~B & ~C &  D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[1184] =  A & ~B & ~C &  D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1185] =  A & ~B & ~C &  D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1186] =  A & ~B & ~C &  D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1187] =  A & ~B & ~C &  D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1188] =  A & ~B & ~C &  D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1189] =  A & ~B & ~C &  D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1190] =  A & ~B & ~C &  D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1191] =  A & ~B & ~C &  D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[1192] =  A & ~B & ~C &  D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1193] =  A & ~B & ~C &  D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1194] =  A & ~B & ~C &  D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1195] =  A & ~B & ~C &  D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[1196] =  A & ~B & ~C &  D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1197] =  A & ~B & ~C &  D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[1198] =  A & ~B & ~C &  D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[1199] =  A & ~B & ~C &  D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[1200] =  A & ~B & ~C &  D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1201] =  A & ~B & ~C &  D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1202] =  A & ~B & ~C &  D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1203] =  A & ~B & ~C &  D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[1204] =  A & ~B & ~C &  D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1205] =  A & ~B & ~C &  D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[1206] =  A & ~B & ~C &  D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[1207] =  A & ~B & ~C &  D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[1208] =  A & ~B & ~C &  D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1209] =  A & ~B & ~C &  D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[1210] =  A & ~B & ~C &  D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[1211] =  A & ~B & ~C &  D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[1212] =  A & ~B & ~C &  D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[1213] =  A & ~B & ~C &  D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[1214] =  A & ~B & ~C &  D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[1215] =  A & ~B & ~C &  D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[1216] =  A & ~B & ~C &  D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1217] =  A & ~B & ~C &  D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1218] =  A & ~B & ~C &  D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1219] =  A & ~B & ~C &  D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1220] =  A & ~B & ~C &  D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1221] =  A & ~B & ~C &  D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1222] =  A & ~B & ~C &  D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1223] =  A & ~B & ~C &  D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1224] =  A & ~B & ~C &  D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1225] =  A & ~B & ~C &  D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1226] =  A & ~B & ~C &  D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1227] =  A & ~B & ~C &  D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1228] =  A & ~B & ~C &  D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1229] =  A & ~B & ~C &  D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1230] =  A & ~B & ~C &  D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1231] =  A & ~B & ~C &  D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[1232] =  A & ~B & ~C &  D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1233] =  A & ~B & ~C &  D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1234] =  A & ~B & ~C &  D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1235] =  A & ~B & ~C &  D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1236] =  A & ~B & ~C &  D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1237] =  A & ~B & ~C &  D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1238] =  A & ~B & ~C &  D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1239] =  A & ~B & ~C &  D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[1240] =  A & ~B & ~C &  D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1241] =  A & ~B & ~C &  D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1242] =  A & ~B & ~C &  D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1243] =  A & ~B & ~C &  D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[1244] =  A & ~B & ~C &  D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1245] =  A & ~B & ~C &  D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[1246] =  A & ~B & ~C &  D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[1247] =  A & ~B & ~C &  D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[1248] =  A & ~B & ~C &  D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1249] =  A & ~B & ~C &  D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1250] =  A & ~B & ~C &  D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1251] =  A & ~B & ~C &  D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1252] =  A & ~B & ~C &  D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1253] =  A & ~B & ~C &  D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1254] =  A & ~B & ~C &  D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1255] =  A & ~B & ~C &  D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[1256] =  A & ~B & ~C &  D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1257] =  A & ~B & ~C &  D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1258] =  A & ~B & ~C &  D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1259] =  A & ~B & ~C &  D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[1260] =  A & ~B & ~C &  D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1261] =  A & ~B & ~C &  D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[1262] =  A & ~B & ~C &  D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[1263] =  A & ~B & ~C &  D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[1264] =  A & ~B & ~C &  D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1265] =  A & ~B & ~C &  D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1266] =  A & ~B & ~C &  D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1267] =  A & ~B & ~C &  D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[1268] =  A & ~B & ~C &  D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1269] =  A & ~B & ~C &  D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[1270] =  A & ~B & ~C &  D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[1271] =  A & ~B & ~C &  D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[1272] =  A & ~B & ~C &  D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1273] =  A & ~B & ~C &  D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[1274] =  A & ~B & ~C &  D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[1275] =  A & ~B & ~C &  D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[1276] =  A & ~B & ~C &  D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[1277] =  A & ~B & ~C &  D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[1278] =  A & ~B & ~C &  D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[1279] =  A & ~B & ~C &  D &  E &  F &  G &  H &  I &  J &  K;
	assign out[1280] =  A & ~B &  C & ~D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1281] =  A & ~B &  C & ~D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1282] =  A & ~B &  C & ~D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1283] =  A & ~B &  C & ~D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1284] =  A & ~B &  C & ~D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1285] =  A & ~B &  C & ~D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1286] =  A & ~B &  C & ~D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1287] =  A & ~B &  C & ~D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1288] =  A & ~B &  C & ~D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1289] =  A & ~B &  C & ~D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1290] =  A & ~B &  C & ~D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1291] =  A & ~B &  C & ~D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1292] =  A & ~B &  C & ~D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1293] =  A & ~B &  C & ~D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1294] =  A & ~B &  C & ~D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1295] =  A & ~B &  C & ~D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[1296] =  A & ~B &  C & ~D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1297] =  A & ~B &  C & ~D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1298] =  A & ~B &  C & ~D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1299] =  A & ~B &  C & ~D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1300] =  A & ~B &  C & ~D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1301] =  A & ~B &  C & ~D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1302] =  A & ~B &  C & ~D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1303] =  A & ~B &  C & ~D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[1304] =  A & ~B &  C & ~D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1305] =  A & ~B &  C & ~D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1306] =  A & ~B &  C & ~D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1307] =  A & ~B &  C & ~D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[1308] =  A & ~B &  C & ~D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1309] =  A & ~B &  C & ~D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[1310] =  A & ~B &  C & ~D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[1311] =  A & ~B &  C & ~D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[1312] =  A & ~B &  C & ~D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1313] =  A & ~B &  C & ~D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1314] =  A & ~B &  C & ~D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1315] =  A & ~B &  C & ~D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1316] =  A & ~B &  C & ~D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1317] =  A & ~B &  C & ~D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1318] =  A & ~B &  C & ~D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1319] =  A & ~B &  C & ~D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[1320] =  A & ~B &  C & ~D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1321] =  A & ~B &  C & ~D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1322] =  A & ~B &  C & ~D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1323] =  A & ~B &  C & ~D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[1324] =  A & ~B &  C & ~D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1325] =  A & ~B &  C & ~D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[1326] =  A & ~B &  C & ~D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[1327] =  A & ~B &  C & ~D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[1328] =  A & ~B &  C & ~D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1329] =  A & ~B &  C & ~D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1330] =  A & ~B &  C & ~D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1331] =  A & ~B &  C & ~D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[1332] =  A & ~B &  C & ~D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1333] =  A & ~B &  C & ~D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[1334] =  A & ~B &  C & ~D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[1335] =  A & ~B &  C & ~D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[1336] =  A & ~B &  C & ~D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1337] =  A & ~B &  C & ~D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[1338] =  A & ~B &  C & ~D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[1339] =  A & ~B &  C & ~D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[1340] =  A & ~B &  C & ~D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[1341] =  A & ~B &  C & ~D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[1342] =  A & ~B &  C & ~D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[1343] =  A & ~B &  C & ~D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[1344] =  A & ~B &  C & ~D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1345] =  A & ~B &  C & ~D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1346] =  A & ~B &  C & ~D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1347] =  A & ~B &  C & ~D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1348] =  A & ~B &  C & ~D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1349] =  A & ~B &  C & ~D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1350] =  A & ~B &  C & ~D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1351] =  A & ~B &  C & ~D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1352] =  A & ~B &  C & ~D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1353] =  A & ~B &  C & ~D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1354] =  A & ~B &  C & ~D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1355] =  A & ~B &  C & ~D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1356] =  A & ~B &  C & ~D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1357] =  A & ~B &  C & ~D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1358] =  A & ~B &  C & ~D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1359] =  A & ~B &  C & ~D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[1360] =  A & ~B &  C & ~D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1361] =  A & ~B &  C & ~D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1362] =  A & ~B &  C & ~D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1363] =  A & ~B &  C & ~D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1364] =  A & ~B &  C & ~D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1365] =  A & ~B &  C & ~D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1366] =  A & ~B &  C & ~D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1367] =  A & ~B &  C & ~D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[1368] =  A & ~B &  C & ~D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1369] =  A & ~B &  C & ~D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1370] =  A & ~B &  C & ~D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1371] =  A & ~B &  C & ~D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[1372] =  A & ~B &  C & ~D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1373] =  A & ~B &  C & ~D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[1374] =  A & ~B &  C & ~D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[1375] =  A & ~B &  C & ~D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[1376] =  A & ~B &  C & ~D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1377] =  A & ~B &  C & ~D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1378] =  A & ~B &  C & ~D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1379] =  A & ~B &  C & ~D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1380] =  A & ~B &  C & ~D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1381] =  A & ~B &  C & ~D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1382] =  A & ~B &  C & ~D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1383] =  A & ~B &  C & ~D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[1384] =  A & ~B &  C & ~D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1385] =  A & ~B &  C & ~D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1386] =  A & ~B &  C & ~D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1387] =  A & ~B &  C & ~D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[1388] =  A & ~B &  C & ~D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1389] =  A & ~B &  C & ~D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[1390] =  A & ~B &  C & ~D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[1391] =  A & ~B &  C & ~D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[1392] =  A & ~B &  C & ~D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1393] =  A & ~B &  C & ~D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1394] =  A & ~B &  C & ~D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1395] =  A & ~B &  C & ~D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[1396] =  A & ~B &  C & ~D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1397] =  A & ~B &  C & ~D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[1398] =  A & ~B &  C & ~D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[1399] =  A & ~B &  C & ~D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[1400] =  A & ~B &  C & ~D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1401] =  A & ~B &  C & ~D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[1402] =  A & ~B &  C & ~D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[1403] =  A & ~B &  C & ~D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[1404] =  A & ~B &  C & ~D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[1405] =  A & ~B &  C & ~D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[1406] =  A & ~B &  C & ~D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[1407] =  A & ~B &  C & ~D &  E &  F &  G &  H &  I &  J &  K;
	assign out[1408] =  A & ~B &  C &  D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1409] =  A & ~B &  C &  D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1410] =  A & ~B &  C &  D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1411] =  A & ~B &  C &  D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1412] =  A & ~B &  C &  D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1413] =  A & ~B &  C &  D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1414] =  A & ~B &  C &  D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1415] =  A & ~B &  C &  D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1416] =  A & ~B &  C &  D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1417] =  A & ~B &  C &  D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1418] =  A & ~B &  C &  D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1419] =  A & ~B &  C &  D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1420] =  A & ~B &  C &  D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1421] =  A & ~B &  C &  D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1422] =  A & ~B &  C &  D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1423] =  A & ~B &  C &  D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[1424] =  A & ~B &  C &  D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1425] =  A & ~B &  C &  D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1426] =  A & ~B &  C &  D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1427] =  A & ~B &  C &  D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1428] =  A & ~B &  C &  D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1429] =  A & ~B &  C &  D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1430] =  A & ~B &  C &  D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1431] =  A & ~B &  C &  D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[1432] =  A & ~B &  C &  D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1433] =  A & ~B &  C &  D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1434] =  A & ~B &  C &  D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1435] =  A & ~B &  C &  D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[1436] =  A & ~B &  C &  D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1437] =  A & ~B &  C &  D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[1438] =  A & ~B &  C &  D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[1439] =  A & ~B &  C &  D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[1440] =  A & ~B &  C &  D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1441] =  A & ~B &  C &  D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1442] =  A & ~B &  C &  D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1443] =  A & ~B &  C &  D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1444] =  A & ~B &  C &  D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1445] =  A & ~B &  C &  D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1446] =  A & ~B &  C &  D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1447] =  A & ~B &  C &  D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[1448] =  A & ~B &  C &  D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1449] =  A & ~B &  C &  D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1450] =  A & ~B &  C &  D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1451] =  A & ~B &  C &  D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[1452] =  A & ~B &  C &  D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1453] =  A & ~B &  C &  D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[1454] =  A & ~B &  C &  D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[1455] =  A & ~B &  C &  D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[1456] =  A & ~B &  C &  D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1457] =  A & ~B &  C &  D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1458] =  A & ~B &  C &  D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1459] =  A & ~B &  C &  D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[1460] =  A & ~B &  C &  D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1461] =  A & ~B &  C &  D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[1462] =  A & ~B &  C &  D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[1463] =  A & ~B &  C &  D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[1464] =  A & ~B &  C &  D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1465] =  A & ~B &  C &  D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[1466] =  A & ~B &  C &  D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[1467] =  A & ~B &  C &  D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[1468] =  A & ~B &  C &  D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[1469] =  A & ~B &  C &  D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[1470] =  A & ~B &  C &  D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[1471] =  A & ~B &  C &  D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[1472] =  A & ~B &  C &  D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1473] =  A & ~B &  C &  D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1474] =  A & ~B &  C &  D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1475] =  A & ~B &  C &  D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1476] =  A & ~B &  C &  D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1477] =  A & ~B &  C &  D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1478] =  A & ~B &  C &  D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1479] =  A & ~B &  C &  D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1480] =  A & ~B &  C &  D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1481] =  A & ~B &  C &  D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1482] =  A & ~B &  C &  D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1483] =  A & ~B &  C &  D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1484] =  A & ~B &  C &  D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1485] =  A & ~B &  C &  D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1486] =  A & ~B &  C &  D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1487] =  A & ~B &  C &  D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[1488] =  A & ~B &  C &  D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1489] =  A & ~B &  C &  D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1490] =  A & ~B &  C &  D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1491] =  A & ~B &  C &  D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1492] =  A & ~B &  C &  D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1493] =  A & ~B &  C &  D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1494] =  A & ~B &  C &  D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1495] =  A & ~B &  C &  D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[1496] =  A & ~B &  C &  D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1497] =  A & ~B &  C &  D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1498] =  A & ~B &  C &  D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1499] =  A & ~B &  C &  D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[1500] =  A & ~B &  C &  D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1501] =  A & ~B &  C &  D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[1502] =  A & ~B &  C &  D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[1503] =  A & ~B &  C &  D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[1504] =  A & ~B &  C &  D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1505] =  A & ~B &  C &  D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1506] =  A & ~B &  C &  D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1507] =  A & ~B &  C &  D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1508] =  A & ~B &  C &  D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1509] =  A & ~B &  C &  D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1510] =  A & ~B &  C &  D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1511] =  A & ~B &  C &  D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[1512] =  A & ~B &  C &  D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1513] =  A & ~B &  C &  D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1514] =  A & ~B &  C &  D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1515] =  A & ~B &  C &  D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[1516] =  A & ~B &  C &  D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1517] =  A & ~B &  C &  D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[1518] =  A & ~B &  C &  D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[1519] =  A & ~B &  C &  D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[1520] =  A & ~B &  C &  D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1521] =  A & ~B &  C &  D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1522] =  A & ~B &  C &  D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1523] =  A & ~B &  C &  D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[1524] =  A & ~B &  C &  D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1525] =  A & ~B &  C &  D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[1526] =  A & ~B &  C &  D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[1527] =  A & ~B &  C &  D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[1528] =  A & ~B &  C &  D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1529] =  A & ~B &  C &  D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[1530] =  A & ~B &  C &  D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[1531] =  A & ~B &  C &  D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[1532] =  A & ~B &  C &  D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[1533] =  A & ~B &  C &  D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[1534] =  A & ~B &  C &  D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[1535] =  A & ~B &  C &  D &  E &  F &  G &  H &  I &  J &  K;
	assign out[1536] =  A &  B & ~C & ~D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1537] =  A &  B & ~C & ~D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1538] =  A &  B & ~C & ~D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1539] =  A &  B & ~C & ~D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1540] =  A &  B & ~C & ~D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1541] =  A &  B & ~C & ~D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1542] =  A &  B & ~C & ~D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1543] =  A &  B & ~C & ~D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1544] =  A &  B & ~C & ~D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1545] =  A &  B & ~C & ~D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1546] =  A &  B & ~C & ~D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1547] =  A &  B & ~C & ~D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1548] =  A &  B & ~C & ~D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1549] =  A &  B & ~C & ~D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1550] =  A &  B & ~C & ~D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1551] =  A &  B & ~C & ~D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[1552] =  A &  B & ~C & ~D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1553] =  A &  B & ~C & ~D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1554] =  A &  B & ~C & ~D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1555] =  A &  B & ~C & ~D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1556] =  A &  B & ~C & ~D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1557] =  A &  B & ~C & ~D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1558] =  A &  B & ~C & ~D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1559] =  A &  B & ~C & ~D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[1560] =  A &  B & ~C & ~D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1561] =  A &  B & ~C & ~D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1562] =  A &  B & ~C & ~D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1563] =  A &  B & ~C & ~D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[1564] =  A &  B & ~C & ~D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1565] =  A &  B & ~C & ~D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[1566] =  A &  B & ~C & ~D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[1567] =  A &  B & ~C & ~D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[1568] =  A &  B & ~C & ~D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1569] =  A &  B & ~C & ~D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1570] =  A &  B & ~C & ~D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1571] =  A &  B & ~C & ~D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1572] =  A &  B & ~C & ~D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1573] =  A &  B & ~C & ~D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1574] =  A &  B & ~C & ~D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1575] =  A &  B & ~C & ~D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[1576] =  A &  B & ~C & ~D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1577] =  A &  B & ~C & ~D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1578] =  A &  B & ~C & ~D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1579] =  A &  B & ~C & ~D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[1580] =  A &  B & ~C & ~D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1581] =  A &  B & ~C & ~D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[1582] =  A &  B & ~C & ~D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[1583] =  A &  B & ~C & ~D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[1584] =  A &  B & ~C & ~D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1585] =  A &  B & ~C & ~D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1586] =  A &  B & ~C & ~D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1587] =  A &  B & ~C & ~D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[1588] =  A &  B & ~C & ~D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1589] =  A &  B & ~C & ~D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[1590] =  A &  B & ~C & ~D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[1591] =  A &  B & ~C & ~D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[1592] =  A &  B & ~C & ~D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1593] =  A &  B & ~C & ~D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[1594] =  A &  B & ~C & ~D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[1595] =  A &  B & ~C & ~D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[1596] =  A &  B & ~C & ~D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[1597] =  A &  B & ~C & ~D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[1598] =  A &  B & ~C & ~D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[1599] =  A &  B & ~C & ~D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[1600] =  A &  B & ~C & ~D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1601] =  A &  B & ~C & ~D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1602] =  A &  B & ~C & ~D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1603] =  A &  B & ~C & ~D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1604] =  A &  B & ~C & ~D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1605] =  A &  B & ~C & ~D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1606] =  A &  B & ~C & ~D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1607] =  A &  B & ~C & ~D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1608] =  A &  B & ~C & ~D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1609] =  A &  B & ~C & ~D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1610] =  A &  B & ~C & ~D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1611] =  A &  B & ~C & ~D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1612] =  A &  B & ~C & ~D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1613] =  A &  B & ~C & ~D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1614] =  A &  B & ~C & ~D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1615] =  A &  B & ~C & ~D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[1616] =  A &  B & ~C & ~D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1617] =  A &  B & ~C & ~D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1618] =  A &  B & ~C & ~D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1619] =  A &  B & ~C & ~D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1620] =  A &  B & ~C & ~D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1621] =  A &  B & ~C & ~D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1622] =  A &  B & ~C & ~D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1623] =  A &  B & ~C & ~D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[1624] =  A &  B & ~C & ~D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1625] =  A &  B & ~C & ~D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1626] =  A &  B & ~C & ~D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1627] =  A &  B & ~C & ~D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[1628] =  A &  B & ~C & ~D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1629] =  A &  B & ~C & ~D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[1630] =  A &  B & ~C & ~D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[1631] =  A &  B & ~C & ~D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[1632] =  A &  B & ~C & ~D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1633] =  A &  B & ~C & ~D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1634] =  A &  B & ~C & ~D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1635] =  A &  B & ~C & ~D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1636] =  A &  B & ~C & ~D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1637] =  A &  B & ~C & ~D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1638] =  A &  B & ~C & ~D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1639] =  A &  B & ~C & ~D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[1640] =  A &  B & ~C & ~D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1641] =  A &  B & ~C & ~D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1642] =  A &  B & ~C & ~D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1643] =  A &  B & ~C & ~D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[1644] =  A &  B & ~C & ~D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1645] =  A &  B & ~C & ~D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[1646] =  A &  B & ~C & ~D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[1647] =  A &  B & ~C & ~D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[1648] =  A &  B & ~C & ~D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1649] =  A &  B & ~C & ~D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1650] =  A &  B & ~C & ~D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1651] =  A &  B & ~C & ~D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[1652] =  A &  B & ~C & ~D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1653] =  A &  B & ~C & ~D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[1654] =  A &  B & ~C & ~D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[1655] =  A &  B & ~C & ~D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[1656] =  A &  B & ~C & ~D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1657] =  A &  B & ~C & ~D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[1658] =  A &  B & ~C & ~D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[1659] =  A &  B & ~C & ~D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[1660] =  A &  B & ~C & ~D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[1661] =  A &  B & ~C & ~D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[1662] =  A &  B & ~C & ~D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[1663] =  A &  B & ~C & ~D &  E &  F &  G &  H &  I &  J &  K;
	assign out[1664] =  A &  B & ~C &  D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1665] =  A &  B & ~C &  D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1666] =  A &  B & ~C &  D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1667] =  A &  B & ~C &  D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1668] =  A &  B & ~C &  D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1669] =  A &  B & ~C &  D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1670] =  A &  B & ~C &  D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1671] =  A &  B & ~C &  D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1672] =  A &  B & ~C &  D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1673] =  A &  B & ~C &  D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1674] =  A &  B & ~C &  D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1675] =  A &  B & ~C &  D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1676] =  A &  B & ~C &  D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1677] =  A &  B & ~C &  D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1678] =  A &  B & ~C &  D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1679] =  A &  B & ~C &  D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[1680] =  A &  B & ~C &  D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1681] =  A &  B & ~C &  D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1682] =  A &  B & ~C &  D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1683] =  A &  B & ~C &  D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1684] =  A &  B & ~C &  D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1685] =  A &  B & ~C &  D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1686] =  A &  B & ~C &  D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1687] =  A &  B & ~C &  D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[1688] =  A &  B & ~C &  D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1689] =  A &  B & ~C &  D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1690] =  A &  B & ~C &  D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1691] =  A &  B & ~C &  D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[1692] =  A &  B & ~C &  D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1693] =  A &  B & ~C &  D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[1694] =  A &  B & ~C &  D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[1695] =  A &  B & ~C &  D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[1696] =  A &  B & ~C &  D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1697] =  A &  B & ~C &  D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1698] =  A &  B & ~C &  D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1699] =  A &  B & ~C &  D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1700] =  A &  B & ~C &  D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1701] =  A &  B & ~C &  D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1702] =  A &  B & ~C &  D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1703] =  A &  B & ~C &  D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[1704] =  A &  B & ~C &  D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1705] =  A &  B & ~C &  D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1706] =  A &  B & ~C &  D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1707] =  A &  B & ~C &  D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[1708] =  A &  B & ~C &  D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1709] =  A &  B & ~C &  D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[1710] =  A &  B & ~C &  D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[1711] =  A &  B & ~C &  D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[1712] =  A &  B & ~C &  D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1713] =  A &  B & ~C &  D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1714] =  A &  B & ~C &  D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1715] =  A &  B & ~C &  D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[1716] =  A &  B & ~C &  D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1717] =  A &  B & ~C &  D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[1718] =  A &  B & ~C &  D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[1719] =  A &  B & ~C &  D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[1720] =  A &  B & ~C &  D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1721] =  A &  B & ~C &  D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[1722] =  A &  B & ~C &  D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[1723] =  A &  B & ~C &  D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[1724] =  A &  B & ~C &  D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[1725] =  A &  B & ~C &  D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[1726] =  A &  B & ~C &  D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[1727] =  A &  B & ~C &  D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[1728] =  A &  B & ~C &  D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1729] =  A &  B & ~C &  D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1730] =  A &  B & ~C &  D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1731] =  A &  B & ~C &  D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1732] =  A &  B & ~C &  D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1733] =  A &  B & ~C &  D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1734] =  A &  B & ~C &  D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1735] =  A &  B & ~C &  D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1736] =  A &  B & ~C &  D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1737] =  A &  B & ~C &  D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1738] =  A &  B & ~C &  D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1739] =  A &  B & ~C &  D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1740] =  A &  B & ~C &  D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1741] =  A &  B & ~C &  D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1742] =  A &  B & ~C &  D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1743] =  A &  B & ~C &  D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[1744] =  A &  B & ~C &  D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1745] =  A &  B & ~C &  D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1746] =  A &  B & ~C &  D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1747] =  A &  B & ~C &  D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1748] =  A &  B & ~C &  D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1749] =  A &  B & ~C &  D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1750] =  A &  B & ~C &  D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1751] =  A &  B & ~C &  D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[1752] =  A &  B & ~C &  D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1753] =  A &  B & ~C &  D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1754] =  A &  B & ~C &  D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1755] =  A &  B & ~C &  D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[1756] =  A &  B & ~C &  D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1757] =  A &  B & ~C &  D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[1758] =  A &  B & ~C &  D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[1759] =  A &  B & ~C &  D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[1760] =  A &  B & ~C &  D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1761] =  A &  B & ~C &  D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1762] =  A &  B & ~C &  D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1763] =  A &  B & ~C &  D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1764] =  A &  B & ~C &  D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1765] =  A &  B & ~C &  D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1766] =  A &  B & ~C &  D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1767] =  A &  B & ~C &  D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[1768] =  A &  B & ~C &  D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1769] =  A &  B & ~C &  D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1770] =  A &  B & ~C &  D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1771] =  A &  B & ~C &  D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[1772] =  A &  B & ~C &  D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1773] =  A &  B & ~C &  D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[1774] =  A &  B & ~C &  D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[1775] =  A &  B & ~C &  D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[1776] =  A &  B & ~C &  D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1777] =  A &  B & ~C &  D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1778] =  A &  B & ~C &  D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1779] =  A &  B & ~C &  D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[1780] =  A &  B & ~C &  D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1781] =  A &  B & ~C &  D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[1782] =  A &  B & ~C &  D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[1783] =  A &  B & ~C &  D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[1784] =  A &  B & ~C &  D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1785] =  A &  B & ~C &  D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[1786] =  A &  B & ~C &  D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[1787] =  A &  B & ~C &  D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[1788] =  A &  B & ~C &  D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[1789] =  A &  B & ~C &  D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[1790] =  A &  B & ~C &  D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[1791] =  A &  B & ~C &  D &  E &  F &  G &  H &  I &  J &  K;
	assign out[1792] =  A &  B &  C & ~D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1793] =  A &  B &  C & ~D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1794] =  A &  B &  C & ~D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1795] =  A &  B &  C & ~D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1796] =  A &  B &  C & ~D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1797] =  A &  B &  C & ~D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1798] =  A &  B &  C & ~D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1799] =  A &  B &  C & ~D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1800] =  A &  B &  C & ~D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1801] =  A &  B &  C & ~D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1802] =  A &  B &  C & ~D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1803] =  A &  B &  C & ~D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1804] =  A &  B &  C & ~D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1805] =  A &  B &  C & ~D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1806] =  A &  B &  C & ~D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1807] =  A &  B &  C & ~D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[1808] =  A &  B &  C & ~D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1809] =  A &  B &  C & ~D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1810] =  A &  B &  C & ~D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1811] =  A &  B &  C & ~D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1812] =  A &  B &  C & ~D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1813] =  A &  B &  C & ~D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1814] =  A &  B &  C & ~D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1815] =  A &  B &  C & ~D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[1816] =  A &  B &  C & ~D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1817] =  A &  B &  C & ~D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1818] =  A &  B &  C & ~D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1819] =  A &  B &  C & ~D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[1820] =  A &  B &  C & ~D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1821] =  A &  B &  C & ~D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[1822] =  A &  B &  C & ~D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[1823] =  A &  B &  C & ~D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[1824] =  A &  B &  C & ~D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1825] =  A &  B &  C & ~D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1826] =  A &  B &  C & ~D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1827] =  A &  B &  C & ~D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1828] =  A &  B &  C & ~D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1829] =  A &  B &  C & ~D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1830] =  A &  B &  C & ~D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1831] =  A &  B &  C & ~D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[1832] =  A &  B &  C & ~D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1833] =  A &  B &  C & ~D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1834] =  A &  B &  C & ~D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1835] =  A &  B &  C & ~D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[1836] =  A &  B &  C & ~D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1837] =  A &  B &  C & ~D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[1838] =  A &  B &  C & ~D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[1839] =  A &  B &  C & ~D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[1840] =  A &  B &  C & ~D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1841] =  A &  B &  C & ~D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1842] =  A &  B &  C & ~D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1843] =  A &  B &  C & ~D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[1844] =  A &  B &  C & ~D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1845] =  A &  B &  C & ~D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[1846] =  A &  B &  C & ~D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[1847] =  A &  B &  C & ~D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[1848] =  A &  B &  C & ~D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1849] =  A &  B &  C & ~D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[1850] =  A &  B &  C & ~D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[1851] =  A &  B &  C & ~D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[1852] =  A &  B &  C & ~D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[1853] =  A &  B &  C & ~D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[1854] =  A &  B &  C & ~D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[1855] =  A &  B &  C & ~D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[1856] =  A &  B &  C & ~D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1857] =  A &  B &  C & ~D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1858] =  A &  B &  C & ~D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1859] =  A &  B &  C & ~D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1860] =  A &  B &  C & ~D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1861] =  A &  B &  C & ~D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1862] =  A &  B &  C & ~D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1863] =  A &  B &  C & ~D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1864] =  A &  B &  C & ~D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1865] =  A &  B &  C & ~D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1866] =  A &  B &  C & ~D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1867] =  A &  B &  C & ~D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1868] =  A &  B &  C & ~D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1869] =  A &  B &  C & ~D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1870] =  A &  B &  C & ~D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1871] =  A &  B &  C & ~D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[1872] =  A &  B &  C & ~D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1873] =  A &  B &  C & ~D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1874] =  A &  B &  C & ~D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1875] =  A &  B &  C & ~D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1876] =  A &  B &  C & ~D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1877] =  A &  B &  C & ~D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1878] =  A &  B &  C & ~D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1879] =  A &  B &  C & ~D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[1880] =  A &  B &  C & ~D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1881] =  A &  B &  C & ~D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1882] =  A &  B &  C & ~D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1883] =  A &  B &  C & ~D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[1884] =  A &  B &  C & ~D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1885] =  A &  B &  C & ~D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[1886] =  A &  B &  C & ~D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[1887] =  A &  B &  C & ~D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[1888] =  A &  B &  C & ~D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1889] =  A &  B &  C & ~D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1890] =  A &  B &  C & ~D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1891] =  A &  B &  C & ~D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1892] =  A &  B &  C & ~D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1893] =  A &  B &  C & ~D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1894] =  A &  B &  C & ~D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1895] =  A &  B &  C & ~D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[1896] =  A &  B &  C & ~D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1897] =  A &  B &  C & ~D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1898] =  A &  B &  C & ~D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1899] =  A &  B &  C & ~D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[1900] =  A &  B &  C & ~D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1901] =  A &  B &  C & ~D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[1902] =  A &  B &  C & ~D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[1903] =  A &  B &  C & ~D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[1904] =  A &  B &  C & ~D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1905] =  A &  B &  C & ~D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1906] =  A &  B &  C & ~D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1907] =  A &  B &  C & ~D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[1908] =  A &  B &  C & ~D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1909] =  A &  B &  C & ~D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[1910] =  A &  B &  C & ~D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[1911] =  A &  B &  C & ~D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[1912] =  A &  B &  C & ~D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1913] =  A &  B &  C & ~D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[1914] =  A &  B &  C & ~D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[1915] =  A &  B &  C & ~D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[1916] =  A &  B &  C & ~D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[1917] =  A &  B &  C & ~D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[1918] =  A &  B &  C & ~D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[1919] =  A &  B &  C & ~D &  E &  F &  G &  H &  I &  J &  K;
	assign out[1920] =  A &  B &  C &  D & ~E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1921] =  A &  B &  C &  D & ~E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1922] =  A &  B &  C &  D & ~E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1923] =  A &  B &  C &  D & ~E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1924] =  A &  B &  C &  D & ~E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1925] =  A &  B &  C &  D & ~E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1926] =  A &  B &  C &  D & ~E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1927] =  A &  B &  C &  D & ~E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1928] =  A &  B &  C &  D & ~E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1929] =  A &  B &  C &  D & ~E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1930] =  A &  B &  C &  D & ~E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1931] =  A &  B &  C &  D & ~E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1932] =  A &  B &  C &  D & ~E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1933] =  A &  B &  C &  D & ~E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1934] =  A &  B &  C &  D & ~E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1935] =  A &  B &  C &  D & ~E & ~F & ~G &  H &  I &  J &  K;
	assign out[1936] =  A &  B &  C &  D & ~E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[1937] =  A &  B &  C &  D & ~E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[1938] =  A &  B &  C &  D & ~E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[1939] =  A &  B &  C &  D & ~E & ~F &  G & ~H & ~I &  J &  K;
	assign out[1940] =  A &  B &  C &  D & ~E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[1941] =  A &  B &  C &  D & ~E & ~F &  G & ~H &  I & ~J &  K;
	assign out[1942] =  A &  B &  C &  D & ~E & ~F &  G & ~H &  I &  J & ~K;
	assign out[1943] =  A &  B &  C &  D & ~E & ~F &  G & ~H &  I &  J &  K;
	assign out[1944] =  A &  B &  C &  D & ~E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[1945] =  A &  B &  C &  D & ~E & ~F &  G &  H & ~I & ~J &  K;
	assign out[1946] =  A &  B &  C &  D & ~E & ~F &  G &  H & ~I &  J & ~K;
	assign out[1947] =  A &  B &  C &  D & ~E & ~F &  G &  H & ~I &  J &  K;
	assign out[1948] =  A &  B &  C &  D & ~E & ~F &  G &  H &  I & ~J & ~K;
	assign out[1949] =  A &  B &  C &  D & ~E & ~F &  G &  H &  I & ~J &  K;
	assign out[1950] =  A &  B &  C &  D & ~E & ~F &  G &  H &  I &  J & ~K;
	assign out[1951] =  A &  B &  C &  D & ~E & ~F &  G &  H &  I &  J &  K;
	assign out[1952] =  A &  B &  C &  D & ~E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[1953] =  A &  B &  C &  D & ~E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[1954] =  A &  B &  C &  D & ~E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[1955] =  A &  B &  C &  D & ~E &  F & ~G & ~H & ~I &  J &  K;
	assign out[1956] =  A &  B &  C &  D & ~E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[1957] =  A &  B &  C &  D & ~E &  F & ~G & ~H &  I & ~J &  K;
	assign out[1958] =  A &  B &  C &  D & ~E &  F & ~G & ~H &  I &  J & ~K;
	assign out[1959] =  A &  B &  C &  D & ~E &  F & ~G & ~H &  I &  J &  K;
	assign out[1960] =  A &  B &  C &  D & ~E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[1961] =  A &  B &  C &  D & ~E &  F & ~G &  H & ~I & ~J &  K;
	assign out[1962] =  A &  B &  C &  D & ~E &  F & ~G &  H & ~I &  J & ~K;
	assign out[1963] =  A &  B &  C &  D & ~E &  F & ~G &  H & ~I &  J &  K;
	assign out[1964] =  A &  B &  C &  D & ~E &  F & ~G &  H &  I & ~J & ~K;
	assign out[1965] =  A &  B &  C &  D & ~E &  F & ~G &  H &  I & ~J &  K;
	assign out[1966] =  A &  B &  C &  D & ~E &  F & ~G &  H &  I &  J & ~K;
	assign out[1967] =  A &  B &  C &  D & ~E &  F & ~G &  H &  I &  J &  K;
	assign out[1968] =  A &  B &  C &  D & ~E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[1969] =  A &  B &  C &  D & ~E &  F &  G & ~H & ~I & ~J &  K;
	assign out[1970] =  A &  B &  C &  D & ~E &  F &  G & ~H & ~I &  J & ~K;
	assign out[1971] =  A &  B &  C &  D & ~E &  F &  G & ~H & ~I &  J &  K;
	assign out[1972] =  A &  B &  C &  D & ~E &  F &  G & ~H &  I & ~J & ~K;
	assign out[1973] =  A &  B &  C &  D & ~E &  F &  G & ~H &  I & ~J &  K;
	assign out[1974] =  A &  B &  C &  D & ~E &  F &  G & ~H &  I &  J & ~K;
	assign out[1975] =  A &  B &  C &  D & ~E &  F &  G & ~H &  I &  J &  K;
	assign out[1976] =  A &  B &  C &  D & ~E &  F &  G &  H & ~I & ~J & ~K;
	assign out[1977] =  A &  B &  C &  D & ~E &  F &  G &  H & ~I & ~J &  K;
	assign out[1978] =  A &  B &  C &  D & ~E &  F &  G &  H & ~I &  J & ~K;
	assign out[1979] =  A &  B &  C &  D & ~E &  F &  G &  H & ~I &  J &  K;
	assign out[1980] =  A &  B &  C &  D & ~E &  F &  G &  H &  I & ~J & ~K;
	assign out[1981] =  A &  B &  C &  D & ~E &  F &  G &  H &  I & ~J &  K;
	assign out[1982] =  A &  B &  C &  D & ~E &  F &  G &  H &  I &  J & ~K;
	assign out[1983] =  A &  B &  C &  D & ~E &  F &  G &  H &  I &  J &  K;
	assign out[1984] =  A &  B &  C &  D &  E & ~F & ~G & ~H & ~I & ~J & ~K;
	assign out[1985] =  A &  B &  C &  D &  E & ~F & ~G & ~H & ~I & ~J &  K;
	assign out[1986] =  A &  B &  C &  D &  E & ~F & ~G & ~H & ~I &  J & ~K;
	assign out[1987] =  A &  B &  C &  D &  E & ~F & ~G & ~H & ~I &  J &  K;
	assign out[1988] =  A &  B &  C &  D &  E & ~F & ~G & ~H &  I & ~J & ~K;
	assign out[1989] =  A &  B &  C &  D &  E & ~F & ~G & ~H &  I & ~J &  K;
	assign out[1990] =  A &  B &  C &  D &  E & ~F & ~G & ~H &  I &  J & ~K;
	assign out[1991] =  A &  B &  C &  D &  E & ~F & ~G & ~H &  I &  J &  K;
	assign out[1992] =  A &  B &  C &  D &  E & ~F & ~G &  H & ~I & ~J & ~K;
	assign out[1993] =  A &  B &  C &  D &  E & ~F & ~G &  H & ~I & ~J &  K;
	assign out[1994] =  A &  B &  C &  D &  E & ~F & ~G &  H & ~I &  J & ~K;
	assign out[1995] =  A &  B &  C &  D &  E & ~F & ~G &  H & ~I &  J &  K;
	assign out[1996] =  A &  B &  C &  D &  E & ~F & ~G &  H &  I & ~J & ~K;
	assign out[1997] =  A &  B &  C &  D &  E & ~F & ~G &  H &  I & ~J &  K;
	assign out[1998] =  A &  B &  C &  D &  E & ~F & ~G &  H &  I &  J & ~K;
	assign out[1999] =  A &  B &  C &  D &  E & ~F & ~G &  H &  I &  J &  K;
	assign out[2000] =  A &  B &  C &  D &  E & ~F &  G & ~H & ~I & ~J & ~K;
	assign out[2001] =  A &  B &  C &  D &  E & ~F &  G & ~H & ~I & ~J &  K;
	assign out[2002] =  A &  B &  C &  D &  E & ~F &  G & ~H & ~I &  J & ~K;
	assign out[2003] =  A &  B &  C &  D &  E & ~F &  G & ~H & ~I &  J &  K;
	assign out[2004] =  A &  B &  C &  D &  E & ~F &  G & ~H &  I & ~J & ~K;
	assign out[2005] =  A &  B &  C &  D &  E & ~F &  G & ~H &  I & ~J &  K;
	assign out[2006] =  A &  B &  C &  D &  E & ~F &  G & ~H &  I &  J & ~K;
	assign out[2007] =  A &  B &  C &  D &  E & ~F &  G & ~H &  I &  J &  K;
	assign out[2008] =  A &  B &  C &  D &  E & ~F &  G &  H & ~I & ~J & ~K;
	assign out[2009] =  A &  B &  C &  D &  E & ~F &  G &  H & ~I & ~J &  K;
	assign out[2010] =  A &  B &  C &  D &  E & ~F &  G &  H & ~I &  J & ~K;
	assign out[2011] =  A &  B &  C &  D &  E & ~F &  G &  H & ~I &  J &  K;
	assign out[2012] =  A &  B &  C &  D &  E & ~F &  G &  H &  I & ~J & ~K;
	assign out[2013] =  A &  B &  C &  D &  E & ~F &  G &  H &  I & ~J &  K;
	assign out[2014] =  A &  B &  C &  D &  E & ~F &  G &  H &  I &  J & ~K;
	assign out[2015] =  A &  B &  C &  D &  E & ~F &  G &  H &  I &  J &  K;
	assign out[2016] =  A &  B &  C &  D &  E &  F & ~G & ~H & ~I & ~J & ~K;
	assign out[2017] =  A &  B &  C &  D &  E &  F & ~G & ~H & ~I & ~J &  K;
	assign out[2018] =  A &  B &  C &  D &  E &  F & ~G & ~H & ~I &  J & ~K;
	assign out[2019] =  A &  B &  C &  D &  E &  F & ~G & ~H & ~I &  J &  K;
	assign out[2020] =  A &  B &  C &  D &  E &  F & ~G & ~H &  I & ~J & ~K;
	assign out[2021] =  A &  B &  C &  D &  E &  F & ~G & ~H &  I & ~J &  K;
	assign out[2022] =  A &  B &  C &  D &  E &  F & ~G & ~H &  I &  J & ~K;
	assign out[2023] =  A &  B &  C &  D &  E &  F & ~G & ~H &  I &  J &  K;
	assign out[2024] =  A &  B &  C &  D &  E &  F & ~G &  H & ~I & ~J & ~K;
	assign out[2025] =  A &  B &  C &  D &  E &  F & ~G &  H & ~I & ~J &  K;
	assign out[2026] =  A &  B &  C &  D &  E &  F & ~G &  H & ~I &  J & ~K;
	assign out[2027] =  A &  B &  C &  D &  E &  F & ~G &  H & ~I &  J &  K;
	assign out[2028] =  A &  B &  C &  D &  E &  F & ~G &  H &  I & ~J & ~K;
	assign out[2029] =  A &  B &  C &  D &  E &  F & ~G &  H &  I & ~J &  K;
	assign out[2030] =  A &  B &  C &  D &  E &  F & ~G &  H &  I &  J & ~K;
	assign out[2031] =  A &  B &  C &  D &  E &  F & ~G &  H &  I &  J &  K;
	assign out[2032] =  A &  B &  C &  D &  E &  F &  G & ~H & ~I & ~J & ~K;
	assign out[2033] =  A &  B &  C &  D &  E &  F &  G & ~H & ~I & ~J &  K;
	assign out[2034] =  A &  B &  C &  D &  E &  F &  G & ~H & ~I &  J & ~K;
	assign out[2035] =  A &  B &  C &  D &  E &  F &  G & ~H & ~I &  J &  K;
	assign out[2036] =  A &  B &  C &  D &  E &  F &  G & ~H &  I & ~J & ~K;
	assign out[2037] =  A &  B &  C &  D &  E &  F &  G & ~H &  I & ~J &  K;
	assign out[2038] =  A &  B &  C &  D &  E &  F &  G & ~H &  I &  J & ~K;
	assign out[2039] =  A &  B &  C &  D &  E &  F &  G & ~H &  I &  J &  K;
	assign out[2040] =  A &  B &  C &  D &  E &  F &  G &  H & ~I & ~J & ~K;
	assign out[2041] =  A &  B &  C &  D &  E &  F &  G &  H & ~I & ~J &  K;
	assign out[2042] =  A &  B &  C &  D &  E &  F &  G &  H & ~I &  J & ~K;
	assign out[2043] =  A &  B &  C &  D &  E &  F &  G &  H & ~I &  J &  K;
	assign out[2044] =  A &  B &  C &  D &  E &  F &  G &  H &  I & ~J & ~K;
	assign out[2045] =  A &  B &  C &  D &  E &  F &  G &  H &  I & ~J &  K;
	assign out[2046] =  A &  B &  C &  D &  E &  F &  G &  H &  I &  J & ~K;
	assign out[2047] =  A &  B &  C &  D &  E &  F &  G &  H &  I &  J &  K;
endmodule